
module fadder (a,b,sub,rm,s); // fadder

