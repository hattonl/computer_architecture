module wallace_tree24 (a, b, z);
    input [23:0]  a, b;
    output [47:0] z;

    
endmodule
